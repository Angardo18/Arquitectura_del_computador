
module divisor(input [31:0] a,b,input clk, output [31:0] q, remainder);

    

end module